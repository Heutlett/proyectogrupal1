module top
(
	// Entradas
	input logic clk_FPGA, reset, start,
	
	// Salidas
	output logic FlagZero, EndFlag, COMFlag, clk_out,
	output logic [7:0] tmp_Serial_ctr,
	output logic [7:0] ReadDataOut
);
	logic clk;
	logic [31:0] WriteData, DataAdr, ReadData;
	logic MemWrite, MemtoReg;
	logic [31:0] PC, Instr;
	
	
	// Clock Manager
	clock_manager clock(
							  .clk_FPGA(clk_FPGA),
							  .reset(reset),
							  .COMFlag(COMFlag),
							  .clk(clk),
							  .tmp_Serial_ctr(tmp_Serial_ctr)
							  );
							  
	// Instancia del procesador
	pipelined_processor cpu(
									// Entradas
									.clk(clk), 
									.reset(reset), 
									.start(start), 
									.Instr(Instr), 
									.ReadData(ReadData), 
									// Salidas
									.MemWrite(MemWrite), 
									.MemtoRegM(MemtoReg),
									.FlagZero(FlagZero),
									.EndFlag(EndFlag),
									.COMFlag(COMFlag),
									.PC(PC), 
									.ALUResult(DataAdr),
									.WriteData(WriteData)
									); 
									
									
	// Memoria de instrucciones
	instr_mem instr_mem(
								// Entradas
								.clk(clk), 
								.InstrAddress(PC),
								// Salidas
								.ReadInstr(Instr)
								);
	
	// Memoria de datos
	data_mem data_mem(
							// Entradas
							.clk(clk), 
							.WriteEnable(MemWrite), 
							.DataAddress(DataAdr), 
							.WriteData(WriteData),
							// Salidas
							.ReadData(ReadData)
							);
	
	interpreter_comunication ic 	(
											// Entradas
											.clk(clk), 
											.reset(reset), 
											.MemtoReg(MemtoReg),
											.COM(COMFlag),
											.ReadData(ReadData),
											// Salidas
											.clk_out(clk_out),
											.ReadDataOut(ReadDataOut)
											);

	
endmodule