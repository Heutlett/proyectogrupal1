package alu_defs;
//--------------------------------------------------------------------
// ALU RESULT TYPES
//--------------------------------------------------------------------
	parameter AND_ =     3'b010;
	parameter OR_ =     	3'b011;
	parameter MOV_ =   	3'b100;
//--------------------------------------------------------------------
// ARITH_UNIT Operations
//--------------------------------------------------------------------
	parameter ARITH_ADD =  3'b000;
	parameter ARITH_SUB =  3'b001;
	parameter ARITH_MUL =  3'b101;
	
endpackage