package alu_defs;
//--------------------------------------------------------------------
// ALU OPERATIONS
//--------------------------------------------------------------------
	
	parameter ARITH_ADD =  	3'b000;
	parameter ARITH_SUB =  	3'b001;
	parameter MOV_ =   		3'b010;
	parameter ARITH_MUL =  	3'b011;
	
endpackage